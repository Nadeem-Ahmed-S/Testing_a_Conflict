module top
  
  initial begin
    $display("Top")
  end
  
endmodule
